`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:16:31 06/26/2016 
// Design Name: 
// Module Name:    receptor_serial 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module receptor_serial(
		input clk,
		input canal_serial,
		
		output reg [7:0] angulo_servo_1,
		output reg [7:0] angulo_servo_2,
		output reg [7:0] angulo_servo_3,
		output reg [7:0] angulo_servo_4
		
    );
	 
	 
	 
	 
	 


endmodule
